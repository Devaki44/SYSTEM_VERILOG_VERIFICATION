# run -all
# 	GENERATOR CLASS DATA
# time=0,data_in=0e,addr=f
# 	DRIVER CLASS DATA
# time=0,data_in=0e,addr=f
# 	MONITOR CLASS DATA
# time=6,clk=1,rst=1,en=1,data_in=0e,addr=f,data_out=00
#     SCOREBOARD CLASS DATA
# time=6,rst=1,en=1,data_in=0e,addr=f,data_out=00
# time=6,rst=1,en=1,data_in=0e,addr=f,out=00
# -----------------------------------------------
# PASS
# -----------------------------------------------
# 	GENERATOR CLASS DATA
# time=6,data_in=07,addr=f
# 	DRIVER CLASS DATA
# time=6,data_in=07,addr=f
# 	MONITOR CLASS DATA
# time=16,clk=1,rst=1,en=0,data_in=07,addr=f,data_out=00
#     SCOREBOARD CLASS DATA
# time=16,rst=1,en=0,data_in=07,addr=f,data_out=00
# time=16,rst=1,en=0,data_in=07,addr=f,out=00
# -----------------------------------------------
# PASS
# -----------------------------------------------
# 	GENERATOR CLASS DATA
# time=16,data_in=11,addr=f
# 	DRIVER CLASS DATA
# time=16,data_in=11,addr=f
# 	MONITOR CLASS DATA
# time=26,clk=1,rst=0,en=1,data_in=11,addr=f,data_out=00
#     SCOREBOARD CLASS DATA
# time=26,rst=0,en=1,data_in=11,addr=f,data_out=00
# time=26,rst=0,en=1,data_in=11,addr=f,out=00
# -----------------------------------------------
# PASS
# -----------------------------------------------
# 	GENERATOR CLASS DATA
# time=26,data_in=00,addr=f
# 	DRIVER CLASS DATA
# time=26,data_in=00,addr=f
# 	MONITOR CLASS DATA
# time=36,clk=1,rst=0,en=0,data_in=00,addr=f,data_out=11
#     SCOREBOARD CLASS DATA
# time=36,rst=0,en=0,data_in=00,addr=f,data_out=11
# time=36,rst=0,en=0,data_in=00,addr=f,out=11
# -----------------------------------------------
# PASS
# -----------------------------------------------
# 	GENERATOR CLASS DATA
# time=36,data_in=09,addr=f
# 	DRIVER CLASS DATA
# time=36,data_in=09,addr=f
# 	MONITOR CLASS DATA
# time=46,clk=1,rst=0,en=1,data_in=09,addr=f,data_out=11
#     SCOREBOARD CLASS DATA
# time=46,rst=0,en=1,data_in=09,addr=f,data_out=11
# time=46,rst=0,en=1,data_in=09,addr=f,out=11
# -----------------------------------------------
# PASS
# -----------------------------------------------
# 	GENERATOR CLASS DATA
# time=46,data_in=0f,addr=f
# 	DRIVER CLASS DATA
# time=46,data_in=0f,addr=f
# 	MONITOR CLASS DATA
# time=56,clk=1,rst=0,en=0,data_in=0f,addr=f,data_out=09
#     SCOREBOARD CLASS DATA
# time=56,rst=0,en=0,data_in=0f,addr=f,data_out=09
# time=56,rst=0,en=0,data_in=0f,addr=f,out=09
# -----------------------------------------------
# PASS
# -----------------------------------------------
# 	GENERATOR CLASS DATA
# time=56,data_in=10,addr=f
# 	DRIVER CLASS DATA
# time=56,data_in=10,addr=f
# 	MONITOR CLASS DATA
# time=66,clk=1,rst=0,en=1,data_in=10,addr=f,data_out=09
#     SCOREBOARD CLASS DATA
# time=66,rst=0,en=1,data_in=10,addr=f,data_out=09
# time=66,rst=0,en=1,data_in=10,addr=f,out=09
# -----------------------------------------------
# PASS
# -----------------------------------------------
# 	GENERATOR CLASS DATA
# time=66,data_in=0c,addr=f
# 	DRIVER CLASS DATA
# time=66,data_in=0c,addr=f
# 	MONITOR CLASS DATA
# time=76,clk=1,rst=0,en=0,data_in=0c,addr=f,data_out=10
#     SCOREBOARD CLASS DATA
# time=76,rst=0,en=0,data_in=0c,addr=f,data_out=10
# time=76,rst=0,en=0,data_in=0c,addr=f,out=10
# -----------------------------------------------
# PASS
# -----------------------------------------------
# 	GENERATOR CLASS DATA
# time=76,data_in=06,addr=f
# 	DRIVER CLASS DATA
# time=76,data_in=06,addr=f
# 	MONITOR CLASS DATA
# time=86,clk=1,rst=0,en=1,data_in=06,addr=f,data_out=10
#     SCOREBOARD CLASS DATA
# time=86,rst=0,en=1,data_in=06,addr=f,data_out=10
# time=86,rst=0,en=1,data_in=06,addr=f,out=10
# -----------------------------------------------
# PASS
# -----------------------------------------------
# 	GENERATOR CLASS DATA
# time=86,data_in=12,addr=f
# 	DRIVER CLASS DATA
# time=86,data_in=12,addr=f
# 	MONITOR CLASS DATA
# time=96,clk=1,rst=0,en=0,data_in=12,addr=f,data_out=06
#     SCOREBOARD CLASS DATA
# time=96,rst=0,en=0,data_in=12,addr=f,data_out=06
# time=96,rst=0,en=0,data_in=12,addr=f,out=06
# -----------------------------------------------
# PASS
# -----------------------------------------------
# 	GENERATOR CLASS DATA
# time=96,data_in=04,addr=f
# 	DRIVER CLASS DATA
# time=96,data_in=04,addr=f
# ** Note: $finish    : testbench.sv(36)
