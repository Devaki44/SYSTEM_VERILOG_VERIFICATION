class transaction;
  bit  clk;
  bit  rst;
  rand bit  t;
  bit  q;
  
endclass
