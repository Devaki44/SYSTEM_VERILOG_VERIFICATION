Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Aug  7 13:03 2025
 GENERATOR CLASS DATA 
time =0,clk=0,rst=1,d=0,q=0
 DRIVER CLASS DATA 
time =5,clk=1,rst=1,d=0,q=0
 MONITOR CLASS DATA 
time =6,clk=1,rst=1,d=0,q=0
 SCOREBOARD CLASS DATA 
time =6,clk=1,rst=1,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =6,clk=1,rst=1,d=1,q=0
 DRIVER CLASS DATA 
time =15,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =16,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =16,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =16,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =25,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =26,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =26,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =26,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =35,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =36,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =36,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =36,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =45,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =46,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =46,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =46,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =55,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =56,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =56,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =56,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =65,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =66,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =66,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =66,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =75,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =76,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =76,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =76,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =85,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =86,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =86,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =86,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =95,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =96,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =96,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =96,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =105,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =106,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =106,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =106,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =115,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =116,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =116,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =116,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =125,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =126,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =126,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =126,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =135,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =136,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =136,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =136,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =145,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =146,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =146,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =146,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =155,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =156,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =156,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =156,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =165,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =166,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =166,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =166,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =175,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =176,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =176,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =176,clk=1,rst=0,d=0,q=0
 DRIVER CLASS DATA 
time =185,clk=1,rst=0,d=0,q=0
 MONITOR CLASS DATA 
time =186,clk=1,rst=0,d=1,q=1
 SCOREBOARD CLASS DATA 
time =186,clk=1,rst=0,d=1,q=1
		PASS		
-----------------------------------------------		
 GENERATOR CLASS DATA 
time =186,clk=1,rst=0,d=1,q=0
 DRIVER CLASS DATA 
time =195,clk=1,rst=0,d=1,q=0
 MONITOR CLASS DATA 
time =196,clk=1,rst=0,d=0,q=0
 SCOREBOARD CLASS DATA 
time =196,clk=1,rst=0,d=0,q=0
		PASS		
-----------------------------------------------		
$finish at simulation time                  196
           V C S   S i m u l a t i o n   R e p o r t 
