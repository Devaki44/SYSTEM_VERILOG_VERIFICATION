interface intf(input logic clk,input logic rst);
  
  logic t;
  logic q;
  
endinterface
