GENERATOR CLASS  
time=0,rst=0,t=0,q=0
  MONITOR CLASS DATA  
time=7,clk=1,rst=1,t=0,q=0
  SCOREBOARD CLASS DATA  
time=7,rst=1,t=0,q=0
time=7,rst=1,t=0,out=0
--------------------------------------------------------------------------------------
PASS
--------------------------------------------------------------------------------------
  GENERATOR CLASS  
time=7,rst=0,t=1,q=0
  DRIVER CLASS  
time=11,clk=0,rst=1,t=1,q=0
  MONITOR CLASS DATA  
time=17,clk=1,rst=1,t=1,q=0
  SCOREBOARD CLASS DATA  
time=17,rst=1,t=1,q=0
time=17,rst=1,t=1,out=0
--------------------------------------------------------------------------------------
PASS
--------------------------------------------------------------------------------------
  GENERATOR CLASS  
time=17,rst=0,t=0,q=0
  DRIVER CLASS  
time=21,clk=0,rst=0,t=0,q=0
  MONITOR CLASS DATA  
time=27,clk=1,rst=0,t=0,q=0
  SCOREBOARD CLASS DATA  
time=27,rst=0,t=0,q=0
time=27,rst=0,t=0,out=0
--------------------------------------------------------------------------------------
PASS
--------------------------------------------------------------------------------------
  GENERATOR CLASS  
time=27,rst=0,t=0,q=0
  DRIVER CLASS  
time=31,clk=0,rst=0,t=0,q=0
  MONITOR CLASS DATA  
time=37,clk=1,rst=0,t=0,q=0
  SCOREBOARD CLASS DATA  
time=37,rst=0,t=0,q=0
time=37,rst=0,t=0,out=0
--------------------------------------------------------------------------------------
PASS
--------------------------------------------------------------------------------------
  GENERATOR CLASS  
time=37,rst=0,t=1,q=0
  DRIVER CLASS  
time=41,clk=0,rst=0,t=1,q=0
  MONITOR CLASS DATA  
time=47,clk=1,rst=0,t=1,q=1
  SCOREBOARD CLASS DATA  
time=47,rst=0,t=1,q=1
time=47,rst=0,t=1,out=1
--------------------------------------------------------------------------------------
PASS
--------------------------------------------------------------------------------------
  GENERATOR CLASS  
time=47,rst=0,t=1,q=0
  DRIVER CLASS  
time=51,clk=0,rst=0,t=1,q=0
  MONITOR CLASS DATA  
time=57,clk=1,rst=0,t=1,q=0
  SCOREBOARD CLASS DATA  
time=57,rst=0,t=1,q=0
time=57,rst=0,t=1,out=0
--------------------------------------------------------------------------------------
PASS
--------------------------------------------------------------------------------------
  GENERATOR CLASS  
time=57,rst=0,t=1,q=0
  DRIVER CLASS  
time=61,clk=0,rst=0,t=1,q=0
  MONITOR CLASS DATA  
time=67,clk=1,rst=0,t=1,q=1
  SCOREBOARD CLASS DATA  
time=67,rst=0,t=1,q=1
time=67,rst=0,t=1,out=1
--------------------------------------------------------------------------------------
PASS
--------------------------------------------------------------------------------------
  GENERATOR CLASS  
time=67,rst=0,t=1,q=0
  DRIVER CLASS  
time=71,clk=0,rst=0,t=1,q=0
  MONITOR CLASS DATA  
time=77,clk=1,rst=0,t=1,q=0
  SCOREBOARD CLASS DATA  
time=77,rst=0,t=1,q=0
time=77,rst=0,t=1,out=0
--------------------------------------------------------------------------------------
PASS
--------------------------------------------------------------------------------------
  GENERATOR CLASS  
time=77,rst=0,t=0,q=0
  DRIVER CLASS  
time=81,clk=0,rst=0,t=0,q=0
  MONITOR CLASS DATA  
time=87,clk=1,rst=0,t=0,q=0
  SCOREBOARD CLASS DATA  
time=87,rst=0,t=0,q=0
time=87,rst=0,t=0,out=0
--------------------------------------------------------------------------------------
PASS
--------------------------------------------------------------------------------------
  GENERATOR CLASS  
time=87,rst=0,t=1,q=0
  DRIVER CLASS  
time=91,clk=0,rst=0,t=1,q=0
  MONITOR CLASS DATA  
time=97,clk=1,rst=0,t=1,q=1
  SCOREBOARD CLASS DATA  
time=97,rst=0,t=1,q=1
time=97,rst=0,t=1,out=1
--------------------------------------------------------------------------------------
PASS
--------------------------------------------------------------------------------------
  GENERATOR CLASS  
time=97,rst=0,t=0,q=0
  DRIVER CLASS  
time=101,clk=0,rst=0,t=0,q=0
  MONITOR CLASS DATA  
time=107,clk=1,rst=0,t=0,q=1
  SCOREBOARD CLASS DATA  
time=107,rst=0,t=0,q=1
time=107,rst=0,t=0,out=1
--------------------------------------------------------------------------------------
PASS
--------------------------------------------------------------------------------------
  GENERATOR CLASS  
time=107,rst=0,t=0,q=0
  DRIVER CLASS  
time=111,clk=0,rst=0,t=0,q=0
  MONITOR CLASS DATA  
time=117,clk=1,rst=0,t=0,q=1
  SCOREBOARD CLASS DATA  
time=117,rst=0,t=0,q=1
time=117,rst=0,t=0,out=1
--------------------------------------------------------------------------------------
PASS
--------------------------------------------------------------------------------------
  GENERATOR CLASS  
time=117,rst=0,t=1,q=0
$finish called from file "testbench.sv", line 24.
$finish at simulation time                  120
           V C S   S i m u l a t i o n   R e p o r t 
