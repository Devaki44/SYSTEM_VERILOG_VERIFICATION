class transaction;
  bit clk;
  bit rst;
  bit en;
  rand bit[3:0] data_in ;
  bit [3:0]data_out;
  bit full;
  bit empty;

endclass
  
