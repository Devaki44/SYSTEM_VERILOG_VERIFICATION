# run -all
#  generator class signals
#  a=1, b=1, c=0, sum =0, carry=0 
#  driver class signals 
#  a=1, b=1, c=0, sum =0, carry=0 
#  monitor class signals 
#  a=1, b=1, c=0, sum =0, carry=1 
#  Scoreboard signals 
#  PASS 
