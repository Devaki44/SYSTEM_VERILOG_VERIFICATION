xcelium> run
 generator class data
time=0, a=1,b=0,sum=0,carry=0
 driver class data
time=0, a=1,b=0,sum=0,carry=0
monitor class data
time=2, a=1,b=0,sum=1,carry=0
 scoreboard class signals
time=2, a=1,b=0,sum=1,carry=0
PASS
 generator class data
time=5, a=0,b=1,sum=0,carry=0
 driver class data
time=5, a=0,b=1,sum=0,carry=0
monitor class data
time=7, a=0,b=1,sum=1,carry=0
 scoreboard class signals
time=7, a=0,b=1,sum=1,carry=0
PASS
Simulation complete via implicit call to $finish(1) at time 12 NS + 1
./test.sv:3 program test(intf vintf);
xcelium> exit
