xcelium> run
  GENERATOR CLASS DATA  
$time = 0,rst = 0,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 0,rst = 0,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 10,clk=0,rst = 1,up_down = 1,count = 0000
  SCOREBOARD CLASS DATA  
$time = 10,rst = 1,up_down = 1,count = 0000
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 10,rst = 0,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 10,rst = 0,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 20,clk=0,rst = 0,up_down = 1,count = 0001
  SCOREBOARD CLASS DATA  
$time = 20,rst = 0,up_down = 1,count = 0001
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 20,rst = 0,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 20,rst = 0,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 30,clk=0,rst = 0,up_down = 1,count = 0010
  SCOREBOARD CLASS DATA  
$time = 30,rst = 0,up_down = 1,count = 0010
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 30,rst = 1,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 30,rst = 1,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 40,clk=0,rst = 1,up_down = 1,count = 0000
  SCOREBOARD CLASS DATA  
$time = 40,rst = 1,up_down = 1,count = 0000
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 40,rst = 0,up_down = 0,count = 0000
  DRIVER CLASS DATA  
$time = 40,rst = 0,up_down = 0,count =0000
  MONITOR CLASS DATA  
$time = 50,clk=0,rst = 0,up_down = 0,count = 1111
  SCOREBOARD CLASS DATA  
$time = 50,rst = 0,up_down = 0,count = 1111
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 50,rst = 1,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 50,rst = 1,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 60,clk=0,rst = 1,up_down = 1,count = 0000
  SCOREBOARD CLASS DATA  
$time = 60,rst = 1,up_down = 1,count = 0000
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 60,rst = 0,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 60,rst = 0,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 70,clk=0,rst = 0,up_down = 1,count = 0001
  SCOREBOARD CLASS DATA  
$time = 70,rst = 0,up_down = 1,count = 0001
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 70,rst = 1,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 70,rst = 1,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 80,clk=0,rst = 1,up_down = 1,count = 0000
  SCOREBOARD CLASS DATA  
$time = 80,rst = 1,up_down = 1,count = 0000
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 80,rst = 0,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 80,rst = 0,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 90,clk=0,rst = 0,up_down = 1,count = 0001
  SCOREBOARD CLASS DATA  
$time = 90,rst = 0,up_down = 1,count = 0001
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 90,rst = 1,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 90,rst = 1,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 100,clk=0,rst = 1,up_down = 1,count = 0000
  SCOREBOARD CLASS DATA  
$time = 100,rst = 1,up_down = 1,count = 0000
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 100,rst = 1,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 100,rst = 1,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 110,clk=0,rst = 1,up_down = 1,count = 0000
  SCOREBOARD CLASS DATA  
$time = 110,rst = 1,up_down = 1,count = 0000
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 110,rst = 0,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 110,rst = 0,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 120,clk=0,rst = 0,up_down = 1,count = 0001
  SCOREBOARD CLASS DATA  
$time = 120,rst = 0,up_down = 1,count = 0001
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 120,rst = 1,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 120,rst = 1,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 130,clk=0,rst = 1,up_down = 1,count = 0000
  SCOREBOARD CLASS DATA  
$time = 130,rst = 1,up_down = 1,count = 0000
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 130,rst = 1,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 130,rst = 1,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 140,clk=0,rst = 1,up_down = 1,count = 0000
  SCOREBOARD CLASS DATA  
$time = 140,rst = 1,up_down = 1,count = 0000
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 140,rst = 1,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 140,rst = 1,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 150,clk=0,rst = 1,up_down = 1,count = 0000
  SCOREBOARD CLASS DATA  
$time = 150,rst = 1,up_down = 1,count = 0000
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 150,rst = 0,up_down = 0,count = 0000
  DRIVER CLASS DATA  
$time = 150,rst = 0,up_down = 0,count =0000
  MONITOR CLASS DATA  
$time = 160,clk=0,rst = 0,up_down = 0,count = 1111
  SCOREBOARD CLASS DATA  
$time = 160,rst = 0,up_down = 0,count = 1111
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 160,rst = 1,up_down = 1,count = 0000
  DRIVER CLASS DATA  
$time = 160,rst = 1,up_down = 1,count =0000
  MONITOR CLASS DATA  
$time = 170,clk=0,rst = 1,up_down = 1,count = 0000
  SCOREBOARD CLASS DATA  
$time = 170,rst = 1,up_down = 1,count = 0000
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 170,rst = 1,up_down = 0,count = 0000
  DRIVER CLASS DATA  
$time = 170,rst = 1,up_down = 0,count =0000
  MONITOR CLASS DATA  
$time = 180,clk=0,rst = 1,up_down = 0,count = 0000
  SCOREBOARD CLASS DATA  
$time = 180,rst = 1,up_down = 0,count = 0000
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 180,rst = 1,up_down = 0,count = 0000
  DRIVER CLASS DATA  
$time = 180,rst = 1,up_down = 0,count =0000
  MONITOR CLASS DATA  
$time = 190,clk=0,rst = 1,up_down = 0,count = 0000
  SCOREBOARD CLASS DATA  
$time = 190,rst = 1,up_down = 0,count = 0000
---------------------PASS--------------------
  GENERATOR CLASS DATA  
$time = 190,rst = 1,up_down = 0,count = 0000
  DRIVER CLASS DATA  
$time = 190,rst = 1,up_down = 0,count =0000
  MONITOR CLASS DATA  
$time = 200,clk=0,rst = 1,up_down = 0,count = 0000
  SCOREBOARD CLASS DATA  
$time = 200,rst = 1,up_down = 0,count = 0000
---------------------PASS--------------------
Simulation complete via implicit call to $finish(1) at time 200 NS + 2
./test.sv:3 program test(intf vintf);
xcelium> exit
