interface intf(input logic clk);

  logic rst;
  logic up_down;
  logic [3:0]count;
endinterface
