interface intf(input logic clk,rst);
  logic d;
  logic q;
endinterface
